`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    13:46:41 05/11/2016
// Design Name:
// Module Name:    font_rom
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module font_rom(
  input [7:0] ascii_i,
  input [3:0] vga_y,
  output reg [7:0] pixels
    );

  always @ ( * ) begin
    case({ascii_i, vga_y})
		12'b00100000_0000: pixels <= 8'b00000000; // 0
		12'b00100000_0001: pixels <= 8'b00000000; // 1
		12'b00100000_0010: pixels <= 8'b00000000; // 2
		12'b00100000_0011: pixels <= 8'b00000000; // 3
		12'b00100000_0100: pixels <= 8'b00000000; // 4
		12'b00100000_0101: pixels <= 8'b00000000; // 5
		12'b00100000_0110: pixels <= 8'b00000000; // 6
		12'b00100000_0111: pixels <= 8'b00000000; // 7
		12'b00100000_1000: pixels <= 8'b00000000; // 8
		12'b00100000_1001: pixels <= 8'b00000000; // 9
		12'b00100000_1010: pixels <= 8'b00000000; // a
		12'b00100000_1011: pixels <= 8'b00000000; // b
		12'b00100000_1100: pixels <= 8'b00000000; // c
		12'b00100000_1101: pixels <= 8'b00000000; // d
		12'b00100000_1110: pixels <= 8'b00000000; // e
		12'b00100000_1111: pixels <= 8'b00000000; // f

		12'b00100010_0000: pixels <= 8'b00000000; // 0
		12'b00100010_0001: pixels <= 8'b01100110; // 1  **  **
		12'b00100010_0010: pixels <= 8'b01100110; // 2  **  **
		12'b00100010_0011: pixels <= 8'b01100110; // 3  **  **
		12'b00100010_0100: pixels <= 8'b00100100; // 4   *  *
		12'b00100010_0101: pixels <= 8'b00000000; // 5
		12'b00100010_0110: pixels <= 8'b00000000; // 6
		12'b00100010_0111: pixels <= 8'b00000000; // 7
		12'b00100010_1000: pixels <= 8'b00000000; // 8
		12'b00100010_1001: pixels <= 8'b00000000; // 9
		12'b00100010_1010: pixels <= 8'b00000000; // a
		12'b00100010_1011: pixels <= 8'b00000000; // b
		12'b00100010_1100: pixels <= 8'b00000000; // c
		12'b00100010_1101: pixels <= 8'b00000000; // d
		12'b00100010_1110: pixels <= 8'b00000000; // e
		12'b00100010_1111: pixels <= 8'b00000000; // f

		12'b00101100_0000: pixels <= 8'b00000000; // 0
		12'b00101100_0001: pixels <= 8'b00000000; // 1
		12'b00101100_0010: pixels <= 8'b00000000; // 2
		12'b00101100_0011: pixels <= 8'b00000000; // 3
		12'b00101100_0100: pixels <= 8'b00000000; // 4
		12'b00101100_0101: pixels <= 8'b00000000; // 5
		12'b00101100_0110: pixels <= 8'b00000000; // 6
		12'b00101100_0111: pixels <= 8'b00000000; // 7
		12'b00101100_1000: pixels <= 8'b00000000; // 8
		12'b00101100_1001: pixels <= 8'b00011000; // 9    **
		12'b00101100_1010: pixels <= 8'b00011000; // a    **
		12'b00101100_1011: pixels <= 8'b00011000; // b    **
		12'b00101100_1100: pixels <= 8'b00110000; // c   **
		12'b00101100_1101: pixels <= 8'b00000000; // d
		12'b00101100_1110: pixels <= 8'b00000000; // e
		12'b00101100_1111: pixels <= 8'b00000000; // f

		12'b00101110_0000: pixels <= 8'b00000000; // 0
		12'b00101110_0001: pixels <= 8'b00000000; // 1
		12'b00101110_0010: pixels <= 8'b00000000; // 2
		12'b00101110_0011: pixels <= 8'b00000000; // 3
		12'b00101110_0100: pixels <= 8'b00000000; // 4
		12'b00101110_0101: pixels <= 8'b00000000; // 5
		12'b00101110_0110: pixels <= 8'b00000000; // 6
		12'b00101110_0111: pixels <= 8'b00000000; // 7
		12'b00101110_1000: pixels <= 8'b00000000; // 8
		12'b00101110_1001: pixels <= 8'b00000000; // 9
		12'b00101110_1010: pixels <= 8'b00011000; // a    **
		12'b00101110_1011: pixels <= 8'b00011000; // b    **
		12'b00101110_1100: pixels <= 8'b00000000; // c
		12'b00101110_1101: pixels <= 8'b00000000; // d
		12'b00101110_1110: pixels <= 8'b00000000; // e
		12'b00101110_1111: pixels <= 8'b00000000; // f

		12'b00111111_0000: pixels <= 8'b00000000; // 0
		12'b00111111_0001: pixels <= 8'b00000000; // 1
		12'b00111111_0010: pixels <= 8'b01111100; // 2  *****
		12'b00111111_0011: pixels <= 8'b11000110; // 3 **   **
		12'b00111111_0100: pixels <= 8'b11000110; // 4 **   **
		12'b00111111_0101: pixels <= 8'b00001100; // 5     **
		12'b00111111_0110: pixels <= 8'b00011000; // 6    **
		12'b00111111_0111: pixels <= 8'b00011000; // 7    **
		12'b00111111_1000: pixels <= 8'b00011000; // 8    **
		12'b00111111_1001: pixels <= 8'b00000000; // 9
		12'b00111111_1010: pixels <= 8'b00011000; // a    **
		12'b00111111_1011: pixels <= 8'b00011000; // b    **
		12'b00111111_1100: pixels <= 8'b00000000; // c
		12'b00111111_1101: pixels <= 8'b00000000; // d
		12'b00111111_1110: pixels <= 8'b00000000; // e
		12'b00111111_1111: pixels <= 8'b00000000; // f

		12'b01000001_0000: pixels <= 8'b00000000; // 0
		12'b01000001_0001: pixels <= 8'b00000000; // 1
		12'b01000001_0010: pixels <= 8'b00010000; // 2    *
		12'b01000001_0011: pixels <= 8'b00111000; // 3   ***
		12'b01000001_0100: pixels <= 8'b01101100; // 4  ** **
		12'b01000001_0101: pixels <= 8'b11000110; // 5 **   **
		12'b01000001_0110: pixels <= 8'b11000110; // 6 **   **
		12'b01000001_0111: pixels <= 8'b11111110; // 7 *******
		12'b01000001_1000: pixels <= 8'b11000110; // 8 **   **
		12'b01000001_1001: pixels <= 8'b11000110; // 9 **   **
		12'b01000001_1010: pixels <= 8'b11000110; // a **   **
		12'b01000001_1011: pixels <= 8'b11000110; // b **   **
		12'b01000001_1100: pixels <= 8'b00000000; // c
		12'b01000001_1101: pixels <= 8'b00000000; // d
		12'b01000001_1110: pixels <= 8'b00000000; // e
		12'b01000001_1111: pixels <= 8'b00000000; // f

		12'b01000010_0000: pixels <= 8'b00000000; // 0
		12'b01000010_0001: pixels <= 8'b00000000; // 1
		12'b01000010_0010: pixels <= 8'b11111100; // 2 ******
		12'b01000010_0011: pixels <= 8'b01100110; // 3  **  **
		12'b01000010_0100: pixels <= 8'b01100110; // 4  **  **
		12'b01000010_0101: pixels <= 8'b01100110; // 5  **  **
		12'b01000010_0110: pixels <= 8'b01111100; // 6  *****
		12'b01000010_0111: pixels <= 8'b01100110; // 7  **  **
		12'b01000010_1000: pixels <= 8'b01100110; // 8  **  **
		12'b01000010_1001: pixels <= 8'b01100110; // 9  **  **
		12'b01000010_1010: pixels <= 8'b01100110; // a  **  **
		12'b01000010_1011: pixels <= 8'b11111100; // b ******
		12'b01000010_1100: pixels <= 8'b00000000; // c
		12'b01000010_1101: pixels <= 8'b00000000; // d
		12'b01000010_1110: pixels <= 8'b00000000; // e
		12'b01000010_1111: pixels <= 8'b00000000; // f

		12'b01000011_0000: pixels <= 8'b00000000; // 0
		12'b01000011_0001: pixels <= 8'b00000000; // 1
		12'b01000011_0010: pixels <= 8'b00111100; // 2   ****
		12'b01000011_0011: pixels <= 8'b01100110; // 3  **  **
		12'b01000011_0100: pixels <= 8'b11000010; // 4 **    *
		12'b01000011_0101: pixels <= 8'b11000000; // 5 **
		12'b01000011_0110: pixels <= 8'b11000000; // 6 **
		12'b01000011_0111: pixels <= 8'b11000000; // 7 **
		12'b01000011_1000: pixels <= 8'b11000000; // 8 **
		12'b01000011_1001: pixels <= 8'b11000010; // 9 **    *
		12'b01000011_1010: pixels <= 8'b01100110; // a  **  **
		12'b01000011_1011: pixels <= 8'b00111100; // b   ****
		12'b01000011_1100: pixels <= 8'b00000000; // c
		12'b01000011_1101: pixels <= 8'b00000000; // d
		12'b01000011_1110: pixels <= 8'b00000000; // e
		12'b01000011_1111: pixels <= 8'b00000000; // f

		12'b01000100_0000: pixels <= 8'b00000000; // 0
		12'b01000100_0001: pixels <= 8'b00000000; // 1
		12'b01000100_0010: pixels <= 8'b11111000; // 2 *****
		12'b01000100_0011: pixels <= 8'b01101100; // 3  ** **
		12'b01000100_0100: pixels <= 8'b01100110; // 4  **  **
		12'b01000100_0101: pixels <= 8'b01100110; // 5  **  **
		12'b01000100_0110: pixels <= 8'b01100110; // 6  **  **
		12'b01000100_0111: pixels <= 8'b01100110; // 7  **  **
		12'b01000100_1000: pixels <= 8'b01100110; // 8  **  **
		12'b01000100_1001: pixels <= 8'b01100110; // 9  **  **
		12'b01000100_1010: pixels <= 8'b01101100; // a  ** **
		12'b01000100_1011: pixels <= 8'b11111000; // b *****
		12'b01000100_1100: pixels <= 8'b00000000; // c
		12'b01000100_1101: pixels <= 8'b00000000; // d
		12'b01000100_1110: pixels <= 8'b00000000; // e
		12'b01000100_1111: pixels <= 8'b00000000; // f

		12'b01000101_0000: pixels <= 8'b00000000; // 0
		12'b01000101_0001: pixels <= 8'b00000000; // 1
		12'b01000101_0010: pixels <= 8'b11111110; // 2 *******
		12'b01000101_0011: pixels <= 8'b01100110; // 3  **  **
		12'b01000101_0100: pixels <= 8'b01100010; // 4  **   *
		12'b01000101_0101: pixels <= 8'b01101000; // 5  ** *
		12'b01000101_0110: pixels <= 8'b01111000; // 6  ****
		12'b01000101_0111: pixels <= 8'b01101000; // 7  ** *
		12'b01000101_1000: pixels <= 8'b01100000; // 8  **
		12'b01000101_1001: pixels <= 8'b01100010; // 9  **   *
		12'b01000101_1010: pixels <= 8'b01100110; // a  **  **
		12'b01000101_1011: pixels <= 8'b11111110; // b *******
		12'b01000101_1100: pixels <= 8'b00000000; // c
		12'b01000101_1101: pixels <= 8'b00000000; // d
		12'b01000101_1110: pixels <= 8'b00000000; // e
		12'b01000101_1111: pixels <= 8'b00000000; // f

		12'b01000110_0000: pixels <= 8'b00000000; // 0
		12'b01000110_0001: pixels <= 8'b00000000; // 1
		12'b01000110_0010: pixels <= 8'b11111110; // 2 *******
		12'b01000110_0011: pixels <= 8'b01100110; // 3  **  **
		12'b01000110_0100: pixels <= 8'b01100010; // 4  **   *
		12'b01000110_0101: pixels <= 8'b01101000; // 5  ** *
		12'b01000110_0110: pixels <= 8'b01111000; // 6  ****
		12'b01000110_0111: pixels <= 8'b01101000; // 7  ** *
		12'b01000110_1000: pixels <= 8'b01100000; // 8  **
		12'b01000110_1001: pixels <= 8'b01100000; // 9  **
		12'b01000110_1010: pixels <= 8'b01100000; // a  **
		12'b01000110_1011: pixels <= 8'b11110000; // b ****
		12'b01000110_1100: pixels <= 8'b00000000; // c
		12'b01000110_1101: pixels <= 8'b00000000; // d
		12'b01000110_1110: pixels <= 8'b00000000; // e
		12'b01000110_1111: pixels <= 8'b00000000; // f

		12'b01000111_0000: pixels <= 8'b00000000; // 0
		12'b01000111_0001: pixels <= 8'b00000000; // 1
		12'b01000111_0010: pixels <= 8'b00111100; // 2   ****
		12'b01000111_0011: pixels <= 8'b01100110; // 3  **  **
		12'b01000111_0100: pixels <= 8'b11000010; // 4 **    *
		12'b01000111_0101: pixels <= 8'b11000000; // 5 **
		12'b01000111_0110: pixels <= 8'b11000000; // 6 **
		12'b01000111_0111: pixels <= 8'b11011110; // 7 ** ****
		12'b01000111_1000: pixels <= 8'b11000110; // 8 **   **
		12'b01000111_1001: pixels <= 8'b11000110; // 9 **   **
		12'b01000111_1010: pixels <= 8'b01100110; // a  **  **
		12'b01000111_1011: pixels <= 8'b00111010; // b   *** *
		12'b01000111_1100: pixels <= 8'b00000000; // c
		12'b01000111_1101: pixels <= 8'b00000000; // d
		12'b01000111_1110: pixels <= 8'b00000000; // e
		12'b01000111_1111: pixels <= 8'b00000000; // f

		12'b01001000_0000: pixels <= 8'b00000000; // 0
		12'b01001000_0001: pixels <= 8'b00000000; // 1
		12'b01001000_0010: pixels <= 8'b11000110; // 2 **   **
		12'b01001000_0011: pixels <= 8'b11000110; // 3 **   **
		12'b01001000_0100: pixels <= 8'b11000110; // 4 **   **
		12'b01001000_0101: pixels <= 8'b11000110; // 5 **   **
		12'b01001000_0110: pixels <= 8'b11111110; // 6 *******
		12'b01001000_0111: pixels <= 8'b11000110; // 7 **   **
		12'b01001000_1000: pixels <= 8'b11000110; // 8 **   **
		12'b01001000_1001: pixels <= 8'b11000110; // 9 **   **
		12'b01001000_1010: pixels <= 8'b11000110; // a **   **
		12'b01001000_1011: pixels <= 8'b11000110; // b **   **
		12'b01001000_1100: pixels <= 8'b00000000; // c
		12'b01001000_1101: pixels <= 8'b00000000; // d
		12'b01001000_1110: pixels <= 8'b00000000; // e
		12'b01001000_1111: pixels <= 8'b00000000; // f

		12'b01001001_0000: pixels <= 8'b00000000; // 0
		12'b01001001_0001: pixels <= 8'b00000000; // 1
		12'b01001001_0010: pixels <= 8'b00111100; // 2   ****
		12'b01001001_0011: pixels <= 8'b00011000; // 3    **
		12'b01001001_0100: pixels <= 8'b00011000; // 4    **
		12'b01001001_0101: pixels <= 8'b00011000; // 5    **
		12'b01001001_0110: pixels <= 8'b00011000; // 6    **
		12'b01001001_0111: pixels <= 8'b00011000; // 7    **
		12'b01001001_1000: pixels <= 8'b00011000; // 8    **
		12'b01001001_1001: pixels <= 8'b00011000; // 9    **
		12'b01001001_1010: pixels <= 8'b00011000; // a    **
		12'b01001001_1011: pixels <= 8'b00111100; // b   ****
		12'b01001001_1100: pixels <= 8'b00000000; // c
		12'b01001001_1101: pixels <= 8'b00000000; // d
		12'b01001001_1110: pixels <= 8'b00000000; // e
		12'b01001001_1111: pixels <= 8'b00000000; // f

		12'b01001010_0000: pixels <= 8'b00000000; // 0
		12'b01001010_0001: pixels <= 8'b00000000; // 1
		12'b01001010_0010: pixels <= 8'b00011110; // 2    ****
		12'b01001010_0011: pixels <= 8'b00001100; // 3     **
		12'b01001010_0100: pixels <= 8'b00001100; // 4     **
		12'b01001010_0101: pixels <= 8'b00001100; // 5     **
		12'b01001010_0110: pixels <= 8'b00001100; // 6     **
		12'b01001010_0111: pixels <= 8'b00001100; // 7     **
		12'b01001010_1000: pixels <= 8'b11001100; // 8 **  **
		12'b01001010_1001: pixels <= 8'b11001100; // 9 **  **
		12'b01001010_1010: pixels <= 8'b11001100; // a **  **
		12'b01001010_1011: pixels <= 8'b01111000; // b  ****
		12'b01001010_1100: pixels <= 8'b00000000; // c
		12'b01001010_1101: pixels <= 8'b00000000; // d
		12'b01001010_1110: pixels <= 8'b00000000; // e
		12'b01001010_1111: pixels <= 8'b00000000; // f

		12'b01001011_0000: pixels <= 8'b00000000; // 0
		12'b01001011_0001: pixels <= 8'b00000000; // 1
		12'b01001011_0010: pixels <= 8'b11100110; // 2 ***  **
		12'b01001011_0011: pixels <= 8'b01100110; // 3  **  **
		12'b01001011_0100: pixels <= 8'b01100110; // 4  **  **
		12'b01001011_0101: pixels <= 8'b01101100; // 5  ** **
		12'b01001011_0110: pixels <= 8'b01111000; // 6  ****
		12'b01001011_0111: pixels <= 8'b01111000; // 7  ****
		12'b01001011_1000: pixels <= 8'b01101100; // 8  ** **
		12'b01001011_1001: pixels <= 8'b01100110; // 9  **  **
		12'b01001011_1010: pixels <= 8'b01100110; // a  **  **
		12'b01001011_1011: pixels <= 8'b11100110; // b ***  **
		12'b01001011_1100: pixels <= 8'b00000000; // c
		12'b01001011_1101: pixels <= 8'b00000000; // d
		12'b01001011_1110: pixels <= 8'b00000000; // e
		12'b01001011_1111: pixels <= 8'b00000000; // f

		12'b01001100_0000: pixels <= 8'b00000000; // 0
		12'b01001100_0001: pixels <= 8'b00000000; // 1
		12'b01001100_0010: pixels <= 8'b11110000; // 2 ****
		12'b01001100_0011: pixels <= 8'b01100000; // 3  **
		12'b01001100_0100: pixels <= 8'b01100000; // 4  **
		12'b01001100_0101: pixels <= 8'b01100000; // 5  **
		12'b01001100_0110: pixels <= 8'b01100000; // 6  **
		12'b01001100_0111: pixels <= 8'b01100000; // 7  **
		12'b01001100_1000: pixels <= 8'b01100000; // 8  **
		12'b01001100_1001: pixels <= 8'b01100010; // 9  **   *
		12'b01001100_1010: pixels <= 8'b01100110; // a  **  **
		12'b01001100_1011: pixels <= 8'b11111110; // b *******
		12'b01001100_1100: pixels <= 8'b00000000; // c
		12'b01001100_1101: pixels <= 8'b00000000; // d
		12'b01001100_1110: pixels <= 8'b00000000; // e
		12'b01001100_1111: pixels <= 8'b00000000; // f

		12'b01001101_0000: pixels <= 8'b00000000; // 0
		12'b01001101_0001: pixels <= 8'b00000000; // 1
		12'b01001101_0010: pixels <= 8'b11000011; // 2 **    **
		12'b01001101_0011: pixels <= 8'b11100111; // 3 ***  ***
		12'b01001101_0100: pixels <= 8'b11111111; // 4 ********
		12'b01001101_0101: pixels <= 8'b11111111; // 5 ********
		12'b01001101_0110: pixels <= 8'b11011011; // 6 ** ** **
		12'b01001101_0111: pixels <= 8'b11000011; // 7 **    **
		12'b01001101_1000: pixels <= 8'b11000011; // 8 **    **
		12'b01001101_1001: pixels <= 8'b11000011; // 9 **    **
		12'b01001101_1010: pixels <= 8'b11000011; // a **    **
		12'b01001101_1011: pixels <= 8'b11000011; // b **    **
		12'b01001101_1100: pixels <= 8'b00000000; // c
		12'b01001101_1101: pixels <= 8'b00000000; // d
		12'b01001101_1110: pixels <= 8'b00000000; // e
		12'b01001101_1111: pixels <= 8'b00000000; // f

		12'b01001110_0000: pixels <= 8'b00000000; // 0
		12'b01001110_0001: pixels <= 8'b00000000; // 1
		12'b01001110_0010: pixels <= 8'b11000110; // 2 **   **
		12'b01001110_0011: pixels <= 8'b11100110; // 3 ***  **
		12'b01001110_0100: pixels <= 8'b11110110; // 4 **** **
		12'b01001110_0101: pixels <= 8'b11111110; // 5 *******
		12'b01001110_0110: pixels <= 8'b11011110; // 6 ** ****
		12'b01001110_0111: pixels <= 8'b11001110; // 7 **  ***
		12'b01001110_1000: pixels <= 8'b11000110; // 8 **   **
		12'b01001110_1001: pixels <= 8'b11000110; // 9 **   **
		12'b01001110_1010: pixels <= 8'b11000110; // a **   **
		12'b01001110_1011: pixels <= 8'b11000110; // b **   **
		12'b01001110_1100: pixels <= 8'b00000000; // c
		12'b01001110_1101: pixels <= 8'b00000000; // d
		12'b01001110_1110: pixels <= 8'b00000000; // e
		12'b01001110_1111: pixels <= 8'b00000000; // f

		12'b01001111_0000: pixels <= 8'b00000000; // 0
		12'b01001111_0001: pixels <= 8'b00000000; // 1
		12'b01001111_0010: pixels <= 8'b01111100; // 2  *****
		12'b01001111_0011: pixels <= 8'b11000110; // 3 **   **
		12'b01001111_0100: pixels <= 8'b11000110; // 4 **   **
		12'b01001111_0101: pixels <= 8'b11000110; // 5 **   **
		12'b01001111_0110: pixels <= 8'b11000110; // 6 **   **
		12'b01001111_0111: pixels <= 8'b11000110; // 7 **   **
		12'b01001111_1000: pixels <= 8'b11000110; // 8 **   **
		12'b01001111_1001: pixels <= 8'b11000110; // 9 **   **
		12'b01001111_1010: pixels <= 8'b11000110; // a **   **
		12'b01001111_1011: pixels <= 8'b01111100; // b  *****
		12'b01001111_1100: pixels <= 8'b00000000; // c
		12'b01001111_1101: pixels <= 8'b00000000; // d
		12'b01001111_1110: pixels <= 8'b00000000; // e
		12'b01001111_1111: pixels <= 8'b00000000; // f

		12'b01010000_0000: pixels <= 8'b00000000; // 0
		12'b01010000_0001: pixels <= 8'b00000000; // 1
		12'b01010000_0010: pixels <= 8'b11111100; // 2 ******
		12'b01010000_0011: pixels <= 8'b01100110; // 3  **  **
		12'b01010000_0100: pixels <= 8'b01100110; // 4  **  **
		12'b01010000_0101: pixels <= 8'b01100110; // 5  **  **
		12'b01010000_0110: pixels <= 8'b01111100; // 6  *****
		12'b01010000_0111: pixels <= 8'b01100000; // 7  **
		12'b01010000_1000: pixels <= 8'b01100000; // 8  **
		12'b01010000_1001: pixels <= 8'b01100000; // 9  **
		12'b01010000_1010: pixels <= 8'b01100000; // a  **
		12'b01010000_1011: pixels <= 8'b11110000; // b ****
		12'b01010000_1100: pixels <= 8'b00000000; // c
		12'b01010000_1101: pixels <= 8'b00000000; // d
		12'b01010000_1110: pixels <= 8'b00000000; // e
		12'b01010000_1111: pixels <= 8'b00000000; // f

		12'b01010001_0000: pixels <= 8'b00000000; // 0
		12'b01010001_0001: pixels <= 8'b00000000; // 1
		12'b01010001_0010: pixels <= 8'b01111100; // 2  *****
		12'b01010001_0011: pixels <= 8'b11000110; // 3 **   **
		12'b01010001_0100: pixels <= 8'b11000110; // 4 **   **
		12'b01010001_0101: pixels <= 8'b11000110; // 5 **   **
		12'b01010001_0110: pixels <= 8'b11000110; // 6 **   **
		12'b01010001_0111: pixels <= 8'b11000110; // 7 **   **
		12'b01010001_1000: pixels <= 8'b11000110; // 8 **   **
		12'b01010001_1001: pixels <= 8'b11010110; // 9 ** * **
		12'b01010001_1010: pixels <= 8'b11011110; // a ** ****
		12'b01010001_1011: pixels <= 8'b01111100; // b  *****
		12'b01010001_1100: pixels <= 8'b00001100; // c     **
		12'b01010001_1101: pixels <= 8'b00001110; // d     ***
		12'b01010001_1110: pixels <= 8'b00000000; // e
		12'b01010001_1111: pixels <= 8'b00000000; // f

		12'b01010010_0000: pixels <= 8'b00000000; // 0
		12'b01010010_0001: pixels <= 8'b00000000; // 1
		12'b01010010_0010: pixels <= 8'b11111100; // 2 ******
		12'b01010010_0011: pixels <= 8'b01100110; // 3  **  **
		12'b01010010_0100: pixels <= 8'b01100110; // 4  **  **
		12'b01010010_0101: pixels <= 8'b01100110; // 5  **  **
		12'b01010010_0110: pixels <= 8'b01111100; // 6  *****
		12'b01010010_0111: pixels <= 8'b01101100; // 7  ** **
		12'b01010010_1000: pixels <= 8'b01100110; // 8  **  **
		12'b01010010_1001: pixels <= 8'b01100110; // 9  **  **
		12'b01010010_1010: pixels <= 8'b01100110; // a  **  **
		12'b01010010_1011: pixels <= 8'b11100110; // b ***  **
		12'b01010010_1100: pixels <= 8'b00000000; // c
		12'b01010010_1101: pixels <= 8'b00000000; // d
		12'b01010010_1110: pixels <= 8'b00000000; // e
		12'b01010010_1111: pixels <= 8'b00000000; // f

		12'b01010011_0000: pixels <= 8'b00000000; // 0
		12'b01010011_0001: pixels <= 8'b00000000; // 1
		12'b01010011_0010: pixels <= 8'b01111100; // 2  *****
		12'b01010011_0011: pixels <= 8'b11000110; // 3 **   **
		12'b01010011_0100: pixels <= 8'b11000110; // 4 **   **
		12'b01010011_0101: pixels <= 8'b01100000; // 5  **
		12'b01010011_0110: pixels <= 8'b00111000; // 6   ***
		12'b01010011_0111: pixels <= 8'b00001100; // 7     **
		12'b01010011_1000: pixels <= 8'b00000110; // 8      **
		12'b01010011_1001: pixels <= 8'b11000110; // 9 **   **
		12'b01010011_1010: pixels <= 8'b11000110; // a **   **
		12'b01010011_1011: pixels <= 8'b01111100; // b  *****
		12'b01010011_1100: pixels <= 8'b00000000; // c
		12'b01010011_1101: pixels <= 8'b00000000; // d
		12'b01010011_1110: pixels <= 8'b00000000; // e
		12'b01010011_1111: pixels <= 8'b00000000; // f

		12'b01010100_0000: pixels <= 8'b00000000; // 0
		12'b01010100_0001: pixels <= 8'b00000000; // 1
		12'b01010100_0010: pixels <= 8'b11111111; // 2 ********
		12'b01010100_0011: pixels <= 8'b11011011; // 3 ** ** **
		12'b01010100_0100: pixels <= 8'b10011001; // 4 *  **  *
		12'b01010100_0101: pixels <= 8'b00011000; // 5    **
		12'b01010100_0110: pixels <= 8'b00011000; // 6    **
		12'b01010100_0111: pixels <= 8'b00011000; // 7    **
		12'b01010100_1000: pixels <= 8'b00011000; // 8    **
		12'b01010100_1001: pixels <= 8'b00011000; // 9    **
		12'b01010100_1010: pixels <= 8'b00011000; // a    **
		12'b01010100_1011: pixels <= 8'b00111100; // b   ****
		12'b01010100_1100: pixels <= 8'b00000000; // c
		12'b01010100_1101: pixels <= 8'b00000000; // d
		12'b01010100_1110: pixels <= 8'b00000000; // e
		12'b01010100_1111: pixels <= 8'b00000000; // f

		12'b01010101_0000: pixels <= 8'b00000000; // 0
		12'b01010101_0001: pixels <= 8'b00000000; // 1
		12'b01010101_0010: pixels <= 8'b11000110; // 2 **   **
		12'b01010101_0011: pixels <= 8'b11000110; // 3 **   **
		12'b01010101_0100: pixels <= 8'b11000110; // 4 **   **
		12'b01010101_0101: pixels <= 8'b11000110; // 5 **   **
		12'b01010101_0110: pixels <= 8'b11000110; // 6 **   **
		12'b01010101_0111: pixels <= 8'b11000110; // 7 **   **
		12'b01010101_1000: pixels <= 8'b11000110; // 8 **   **
		12'b01010101_1001: pixels <= 8'b11000110; // 9 **   **
		12'b01010101_1010: pixels <= 8'b11000110; // a **   **
		12'b01010101_1011: pixels <= 8'b01111100; // b  *****
		12'b01010101_1100: pixels <= 8'b00000000; // c
		12'b01010101_1101: pixels <= 8'b00000000; // d
		12'b01010101_1110: pixels <= 8'b00000000; // e
		12'b01010101_1111: pixels <= 8'b00000000; // f

		12'b01010110_0000: pixels <= 8'b00000000; // 0
		12'b01010110_0001: pixels <= 8'b00000000; // 1
		12'b01010110_0010: pixels <= 8'b11000011; // 2 **    **
		12'b01010110_0011: pixels <= 8'b11000011; // 3 **    **
		12'b01010110_0100: pixels <= 8'b11000011; // 4 **    **
		12'b01010110_0101: pixels <= 8'b11000011; // 5 **    **
		12'b01010110_0110: pixels <= 8'b11000011; // 6 **    **
		12'b01010110_0111: pixels <= 8'b11000011; // 7 **    **
		12'b01010110_1000: pixels <= 8'b11000011; // 8 **    **
		12'b01010110_1001: pixels <= 8'b01100110; // 9  **  **
		12'b01010110_1010: pixels <= 8'b00111100; // a   ****
		12'b01010110_1011: pixels <= 8'b00011000; // b    **
		12'b01010110_1100: pixels <= 8'b00000000; // c
		12'b01010110_1101: pixels <= 8'b00000000; // d
		12'b01010110_1110: pixels <= 8'b00000000; // e
		12'b01010110_1111: pixels <= 8'b00000000; // f

		12'b01010111_0000: pixels <= 8'b00000000; // 0
		12'b01010111_0001: pixels <= 8'b00000000; // 1
		12'b01010111_0010: pixels <= 8'b11000011; // 2 **    **
		12'b01010111_0011: pixels <= 8'b11000011; // 3 **    **
		12'b01010111_0100: pixels <= 8'b11000011; // 4 **    **
		12'b01010111_0101: pixels <= 8'b11000011; // 5 **    **
		12'b01010111_0110: pixels <= 8'b11000011; // 6 **    **
		12'b01010111_0111: pixels <= 8'b11011011; // 7 ** ** **
		12'b01010111_1000: pixels <= 8'b11011011; // 8 ** ** **
		12'b01010111_1001: pixels <= 8'b11111111; // 9 ********
		12'b01010111_1010: pixels <= 8'b01100110; // a  **  **
		12'b01010111_1011: pixels <= 8'b01100110; // b  **  **
		12'b01010111_1100: pixels <= 8'b00000000; // c
		12'b01010111_1101: pixels <= 8'b00000000; // d
		12'b01010111_1110: pixels <= 8'b00000000; // e
		12'b01010111_1111: pixels <= 8'b00000000; // f

		12'b01011000_0000: pixels <= 8'b00000000; // 0
		12'b01011000_0001: pixels <= 8'b00000000; // 1
		12'b01011000_0010: pixels <= 8'b11000011; // 2 **    **
		12'b01011000_0011: pixels <= 8'b11000011; // 3 **    **
		12'b01011000_0100: pixels <= 8'b01100110; // 4  **  **
		12'b01011000_0101: pixels <= 8'b00111100; // 5   ****
		12'b01011000_0110: pixels <= 8'b00011000; // 6    **
		12'b01011000_0111: pixels <= 8'b00011000; // 7    **
		12'b01011000_1000: pixels <= 8'b00111100; // 8   ****
		12'b01011000_1001: pixels <= 8'b01100110; // 9  **  **
		12'b01011000_1010: pixels <= 8'b11000011; // a **    **
		12'b01011000_1011: pixels <= 8'b11000011; // b **    **
		12'b01011000_1100: pixels <= 8'b00000000; // c
		12'b01011000_1101: pixels <= 8'b00000000; // d
		12'b01011000_1110: pixels <= 8'b00000000; // e
		12'b01011000_1111: pixels <= 8'b00000000; // f

		12'b01011001_0000: pixels <= 8'b00000000; // 0
		12'b01011001_0001: pixels <= 8'b00000000; // 1
		12'b01011001_0010: pixels <= 8'b11000011; // 2 **    **
		12'b01011001_0011: pixels <= 8'b11000011; // 3 **    **
		12'b01011001_0100: pixels <= 8'b11000011; // 4 **    **
		12'b01011001_0101: pixels <= 8'b01100110; // 5  **  **
		12'b01011001_0110: pixels <= 8'b00111100; // 6   ****
		12'b01011001_0111: pixels <= 8'b00011000; // 7    **
		12'b01011001_1000: pixels <= 8'b00011000; // 8    **
		12'b01011001_1001: pixels <= 8'b00011000; // 9    **
		12'b01011001_1010: pixels <= 8'b00011000; // a    **
		12'b01011001_1011: pixels <= 8'b00111100; // b   ****
		12'b01011001_1100: pixels <= 8'b00000000; // c
		12'b01011001_1101: pixels <= 8'b00000000; // d
		12'b01011001_1110: pixels <= 8'b00000000; // e
		12'b01011001_1111: pixels <= 8'b00000000; // f

		12'b01011010_0000: pixels <= 8'b00000000; // 0
		12'b01011010_0001: pixels <= 8'b00000000; // 1
		12'b01011010_0010: pixels <= 8'b11111111; // 2 ********
		12'b01011010_0011: pixels <= 8'b11000011; // 3 **    **
		12'b01011010_0100: pixels <= 8'b10000110; // 4 *    **
		12'b01011010_0101: pixels <= 8'b00001100; // 5     **
		12'b01011010_0110: pixels <= 8'b00011000; // 6    **
		12'b01011010_0111: pixels <= 8'b00110000; // 7   **
		12'b01011010_1000: pixels <= 8'b01100000; // 8  **
		12'b01011010_1001: pixels <= 8'b11000001; // 9 **     *
		12'b01011010_1010: pixels <= 8'b11000011; // a **    **
		12'b01011010_1011: pixels <= 8'b11111111; // b ********
		12'b01011010_1100: pixels <= 8'b00000000; // c
		12'b01011010_1101: pixels <= 8'b00000000; // d
		12'b01011010_1110: pixels <= 8'b00000000; // e
		12'b01011010_1111: pixels <= 8'b00000000; // f

		12'b01100001_0000: pixels <= 8'b00000000; // 0
		12'b01100001_0001: pixels <= 8'b00000000; // 1
		12'b01100001_0010: pixels <= 8'b00000000; // 2
		12'b01100001_0011: pixels <= 8'b00000000; // 3
		12'b01100001_0100: pixels <= 8'b00000000; // 4
		12'b01100001_0101: pixels <= 8'b01111000; // 5  ****
		12'b01100001_0110: pixels <= 8'b00001100; // 6     **
		12'b01100001_0111: pixels <= 8'b01111100; // 7  *****
		12'b01100001_1000: pixels <= 8'b11001100; // 8 **  **
		12'b01100001_1001: pixels <= 8'b11001100; // 9 **  **
		12'b01100001_1010: pixels <= 8'b11001100; // a **  **
		12'b01100001_1011: pixels <= 8'b01110110; // b  *** **
		12'b01100001_1100: pixels <= 8'b00000000; // c
		12'b01100001_1101: pixels <= 8'b00000000; // d
		12'b01100001_1110: pixels <= 8'b00000000; // e
		12'b01100001_1111: pixels <= 8'b00000000; // f

		12'b01100010_0000: pixels <= 8'b00000000; // 0
		12'b01100010_0001: pixels <= 8'b00000000; // 1
		12'b01100010_0010: pixels <= 8'b11100000; // 2  ***
		12'b01100010_0011: pixels <= 8'b01100000; // 3   **
		12'b01100010_0100: pixels <= 8'b01100000; // 4   **
		12'b01100010_0101: pixels <= 8'b01111000; // 5   ****
		12'b01100010_0110: pixels <= 8'b01101100; // 6   ** **
		12'b01100010_0111: pixels <= 8'b01100110; // 7   **  **
		12'b01100010_1000: pixels <= 8'b01100110; // 8   **  **
		12'b01100010_1001: pixels <= 8'b01100110; // 9   **  **
		12'b01100010_1010: pixels <= 8'b01100110; // a   **  **
		12'b01100010_1011: pixels <= 8'b01111100; // b   *****
		12'b01100010_1100: pixels <= 8'b00000000; // c
		12'b01100010_1101: pixels <= 8'b00000000; // d
		12'b01100010_1110: pixels <= 8'b00000000; // e
		12'b01100010_1111: pixels <= 8'b00000000; // f

		12'b01100011_0000: pixels <= 8'b00000000; // 0
		12'b01100011_0001: pixels <= 8'b00000000; // 1
		12'b01100011_0010: pixels <= 8'b00000000; // 2
		12'b01100011_0011: pixels <= 8'b00000000; // 3
		12'b01100011_0100: pixels <= 8'b00000000; // 4
		12'b01100011_0101: pixels <= 8'b01111100; // 5  *****
		12'b01100011_0110: pixels <= 8'b11000110; // 6 **   **
		12'b01100011_0111: pixels <= 8'b11000000; // 7 **
		12'b01100011_1000: pixels <= 8'b11000000; // 8 **
		12'b01100011_1001: pixels <= 8'b11000000; // 9 **
		12'b01100011_1010: pixels <= 8'b11000110; // a **   **
		12'b01100011_1011: pixels <= 8'b01111100; // b  *****
		12'b01100011_1100: pixels <= 8'b00000000; // c
		12'b01100011_1101: pixels <= 8'b00000000; // d
		12'b01100011_1110: pixels <= 8'b00000000; // e
		12'b01100011_1111: pixels <= 8'b00000000; // f

		12'b01100100_0000: pixels <= 8'b00000000; // 0
		12'b01100100_0001: pixels <= 8'b00000000; // 1
		12'b01100100_0010: pixels <= 8'b00011100; // 2    ***
		12'b01100100_0011: pixels <= 8'b00001100; // 3     **
		12'b01100100_0100: pixels <= 8'b00001100; // 4     **
		12'b01100100_0101: pixels <= 8'b00111100; // 5   ****
		12'b01100100_0110: pixels <= 8'b01101100; // 6  ** **
		12'b01100100_0111: pixels <= 8'b11001100; // 7 **  **
		12'b01100100_1000: pixels <= 8'b11001100; // 8 **  **
		12'b01100100_1001: pixels <= 8'b11001100; // 9 **  **
		12'b01100100_1010: pixels <= 8'b11001100; // a **  **
		12'b01100100_1011: pixels <= 8'b01110110; // b  *** **
		12'b01100100_1100: pixels <= 8'b00000000; // c
		12'b01100100_1101: pixels <= 8'b00000000; // d
		12'b01100100_1110: pixels <= 8'b00000000; // e
		12'b01100100_1111: pixels <= 8'b00000000; // f

		12'b01100101_0000: pixels <= 8'b00000000; // 0
		12'b01100101_0001: pixels <= 8'b00000000; // 1
		12'b01100101_0010: pixels <= 8'b00000000; // 2
		12'b01100101_0011: pixels <= 8'b00000000; // 3
		12'b01100101_0100: pixels <= 8'b00000000; // 4
		12'b01100101_0101: pixels <= 8'b01111100; // 5  *****
		12'b01100101_0110: pixels <= 8'b11000110; // 6 **   **
		12'b01100101_0111: pixels <= 8'b11111110; // 7 *******
		12'b01100101_1000: pixels <= 8'b11000000; // 8 **
		12'b01100101_1001: pixels <= 8'b11000000; // 9 **
		12'b01100101_1010: pixels <= 8'b11000110; // a **   **
		12'b01100101_1011: pixels <= 8'b01111100; // b  *****
		12'b01100101_1100: pixels <= 8'b00000000; // c
		12'b01100101_1101: pixels <= 8'b00000000; // d
		12'b01100101_1110: pixels <= 8'b00000000; // e
		12'b01100101_1111: pixels <= 8'b00000000; // f

		12'b01100110_0000: pixels <= 8'b00000000; // 0
		12'b01100110_0001: pixels <= 8'b00000000; // 1
		12'b01100110_0010: pixels <= 8'b00111000; // 2   ***
		12'b01100110_0011: pixels <= 8'b01101100; // 3  ** **
		12'b01100110_0100: pixels <= 8'b01100100; // 4  **  *
		12'b01100110_0101: pixels <= 8'b01100000; // 5  **
		12'b01100110_0110: pixels <= 8'b11110000; // 6 ****
		12'b01100110_0111: pixels <= 8'b01100000; // 7  **
		12'b01100110_1000: pixels <= 8'b01100000; // 8  **
		12'b01100110_1001: pixels <= 8'b01100000; // 9  **
		12'b01100110_1010: pixels <= 8'b01100000; // a  **
		12'b01100110_1011: pixels <= 8'b11110000; // b ****
		12'b01100110_1100: pixels <= 8'b00000000; // c
		12'b01100110_1101: pixels <= 8'b00000000; // d
		12'b01100110_1110: pixels <= 8'b00000000; // e
		12'b01100110_1111: pixels <= 8'b00000000; // f

		12'b01100111_0000: pixels <= 8'b00000000; // 0
		12'b01100111_0001: pixels <= 8'b00000000; // 1
		12'b01100111_0010: pixels <= 8'b00000000; // 2
		12'b01100111_0011: pixels <= 8'b00000000; // 3
		12'b01100111_0100: pixels <= 8'b00000000; // 4
		12'b01100111_0101: pixels <= 8'b01110110; // 5  *** **
		12'b01100111_0110: pixels <= 8'b11001100; // 6 **  **
		12'b01100111_0111: pixels <= 8'b11001100; // 7 **  **
		12'b01100111_1000: pixels <= 8'b11001100; // 8 **  **
		12'b01100111_1001: pixels <= 8'b11001100; // 9 **  **
		12'b01100111_1010: pixels <= 8'b11001100; // a **  **
		12'b01100111_1011: pixels <= 8'b01111100; // b  *****
		12'b01100111_1100: pixels <= 8'b00001100; // c     **
		12'b01100111_1101: pixels <= 8'b11001100; // d **  **
		12'b01100111_1110: pixels <= 8'b01111000; // e  ****
		12'b01100111_1111: pixels <= 8'b00000000; // f

		12'b01101000_0000: pixels <= 8'b00000000; // 0
		12'b01101000_0001: pixels <= 8'b00000000; // 1
		12'b01101000_0010: pixels <= 8'b11100000; // 2 ***
		12'b01101000_0011: pixels <= 8'b01100000; // 3  **
		12'b01101000_0100: pixels <= 8'b01100000; // 4  **
		12'b01101000_0101: pixels <= 8'b01101100; // 5  ** **
		12'b01101000_0110: pixels <= 8'b01110110; // 6  *** **
		12'b01101000_0111: pixels <= 8'b01100110; // 7  **  **
		12'b01101000_1000: pixels <= 8'b01100110; // 8  **  **
		12'b01101000_1001: pixels <= 8'b01100110; // 9  **  **
		12'b01101000_1010: pixels <= 8'b01100110; // a  **  **
		12'b01101000_1011: pixels <= 8'b11100110; // b ***  **
		12'b01101000_1100: pixels <= 8'b00000000; // c
		12'b01101000_1101: pixels <= 8'b00000000; // d
		12'b01101000_1110: pixels <= 8'b00000000; // e
		12'b01101000_1111: pixels <= 8'b00000000; // f

		12'b01101001_0000: pixels <= 8'b00000000; // 0
		12'b01101001_0001: pixels <= 8'b00000000; // 1
		12'b01101001_0010: pixels <= 8'b00011000; // 2    **
		12'b01101001_0011: pixels <= 8'b00011000; // 3    **
		12'b01101001_0100: pixels <= 8'b00000000; // 4
		12'b01101001_0101: pixels <= 8'b00111000; // 5   ***
		12'b01101001_0110: pixels <= 8'b00011000; // 6    **
		12'b01101001_0111: pixels <= 8'b00011000; // 7    **
		12'b01101001_1000: pixels <= 8'b00011000; // 8    **
		12'b01101001_1001: pixels <= 8'b00011000; // 9    **
		12'b01101001_1010: pixels <= 8'b00011000; // a    **
		12'b01101001_1011: pixels <= 8'b00111100; // b   ****
		12'b01101001_1100: pixels <= 8'b00000000; // c
		12'b01101001_1101: pixels <= 8'b00000000; // d
		12'b01101001_1110: pixels <= 8'b00000000; // e
		12'b01101001_1111: pixels <= 8'b00000000; // f

		12'b01101010_0000: pixels <= 8'b00000000; // 0
		12'b01101010_0001: pixels <= 8'b00000000; // 1
		12'b01101010_0010: pixels <= 8'b00000110; // 2      **
		12'b01101010_0011: pixels <= 8'b00000110; // 3      **
		12'b01101010_0100: pixels <= 8'b00000000; // 4
		12'b01101010_0101: pixels <= 8'b00001110; // 5     ***
		12'b01101010_0110: pixels <= 8'b00000110; // 6      **
		12'b01101010_0111: pixels <= 8'b00000110; // 7      **
		12'b01101010_1000: pixels <= 8'b00000110; // 8      **
		12'b01101010_1001: pixels <= 8'b00000110; // 9      **
		12'b01101010_1010: pixels <= 8'b00000110; // a      **
		12'b01101010_1011: pixels <= 8'b00000110; // b      **
		12'b01101010_1100: pixels <= 8'b01100110; // c  **  **
		12'b01101010_1101: pixels <= 8'b01100110; // d  **  **
		12'b01101010_1110: pixels <= 8'b00111100; // e   ****
		12'b01101010_1111: pixels <= 8'b00000000; // f

		12'b01101011_0000: pixels <= 8'b00000000; // 0
		12'b01101011_0001: pixels <= 8'b00000000; // 1
		12'b01101011_0010: pixels <= 8'b11100000; // 2 ***
		12'b01101011_0011: pixels <= 8'b01100000; // 3  **
		12'b01101011_0100: pixels <= 8'b01100000; // 4  **
		12'b01101011_0101: pixels <= 8'b01100110; // 5  **  **
		12'b01101011_0110: pixels <= 8'b01101100; // 6  ** **
		12'b01101011_0111: pixels <= 8'b01111000; // 7  ****
		12'b01101011_1000: pixels <= 8'b01111000; // 8  ****
		12'b01101011_1001: pixels <= 8'b01101100; // 9  ** **
		12'b01101011_1010: pixels <= 8'b01100110; // a  **  **
		12'b01101011_1011: pixels <= 8'b11100110; // b ***  **
		12'b01101011_1100: pixels <= 8'b00000000; // c
		12'b01101011_1101: pixels <= 8'b00000000; // d
		12'b01101011_1110: pixels <= 8'b00000000; // e
		12'b01101011_1111: pixels <= 8'b00000000; // f

		12'b01101100_0000: pixels <= 8'b00000000; // 0
		12'b01101100_0001: pixels <= 8'b00000000; // 1
		12'b01101100_0010: pixels <= 8'b00111000; // 2   ***
		12'b01101100_0011: pixels <= 8'b00011000; // 3    **
		12'b01101100_0100: pixels <= 8'b00011000; // 4    **
		12'b01101100_0101: pixels <= 8'b00011000; // 5    **
		12'b01101100_0110: pixels <= 8'b00011000; // 6    **
		12'b01101100_0111: pixels <= 8'b00011000; // 7    **
		12'b01101100_1000: pixels <= 8'b00011000; // 8    **
		12'b01101100_1001: pixels <= 8'b00011000; // 9    **
		12'b01101100_1010: pixels <= 8'b00011000; // a    **
		12'b01101100_1011: pixels <= 8'b00111100; // b   ****
		12'b01101100_1100: pixels <= 8'b00000000; // c
		12'b01101100_1101: pixels <= 8'b00000000; // d
		12'b01101100_1110: pixels <= 8'b00000000; // e
		12'b01101100_1111: pixels <= 8'b00000000; // f

		12'b01101101_0000: pixels <= 8'b00000000; // 0
		12'b01101101_0001: pixels <= 8'b00000000; // 1
		12'b01101101_0010: pixels <= 8'b00000000; // 2
		12'b01101101_0011: pixels <= 8'b00000000; // 3
		12'b01101101_0100: pixels <= 8'b00000000; // 4
		12'b01101101_0101: pixels <= 8'b11100110; // 5 ***  **
		12'b01101101_0110: pixels <= 8'b11111111; // 6 ********
		12'b01101101_0111: pixels <= 8'b11011011; // 7 ** ** **
		12'b01101101_1000: pixels <= 8'b11011011; // 8 ** ** **
		12'b01101101_1001: pixels <= 8'b11011011; // 9 ** ** **
		12'b01101101_1010: pixels <= 8'b11011011; // a ** ** **
		12'b01101101_1011: pixels <= 8'b11011011; // b ** ** **
		12'b01101101_1100: pixels <= 8'b00000000; // c
		12'b01101101_1101: pixels <= 8'b00000000; // d
		12'b01101101_1110: pixels <= 8'b00000000; // e
		12'b01101101_1111: pixels <= 8'b00000000; // f

		12'b01101110_0000: pixels <= 8'b00000000; // 0
		12'b01101110_0001: pixels <= 8'b00000000; // 1
		12'b01101110_0010: pixels <= 8'b00000000; // 2
		12'b01101110_0011: pixels <= 8'b00000000; // 3
		12'b01101110_0100: pixels <= 8'b00000000; // 4
		12'b01101110_0101: pixels <= 8'b11011100; // 5 ** ***
		12'b01101110_0110: pixels <= 8'b01100110; // 6  **  **
		12'b01101110_0111: pixels <= 8'b01100110; // 7  **  **
		12'b01101110_1000: pixels <= 8'b01100110; // 8  **  **
		12'b01101110_1001: pixels <= 8'b01100110; // 9  **  **
		12'b01101110_1010: pixels <= 8'b01100110; // a  **  **
		12'b01101110_1011: pixels <= 8'b01100110; // b  **  **
		12'b01101110_1100: pixels <= 8'b00000000; // c
		12'b01101110_1101: pixels <= 8'b00000000; // d
		12'b01101110_1110: pixels <= 8'b00000000; // e
		12'b01101110_1111: pixels <= 8'b00000000; // f

		12'b01101111_0000: pixels <= 8'b00000000; // 0
		12'b01101111_0001: pixels <= 8'b00000000; // 1
		12'b01101111_0010: pixels <= 8'b00000000; // 2
		12'b01101111_0011: pixels <= 8'b00000000; // 3
		12'b01101111_0100: pixels <= 8'b00000000; // 4
		12'b01101111_0101: pixels <= 8'b01111100; // 5  *****
		12'b01101111_0110: pixels <= 8'b11000110; // 6 **   **
		12'b01101111_0111: pixels <= 8'b11000110; // 7 **   **
		12'b01101111_1000: pixels <= 8'b11000110; // 8 **   **
		12'b01101111_1001: pixels <= 8'b11000110; // 9 **   **
		12'b01101111_1010: pixels <= 8'b11000110; // a **   **
		12'b01101111_1011: pixels <= 8'b01111100; // b  *****
		12'b01101111_1100: pixels <= 8'b00000000; // c
		12'b01101111_1101: pixels <= 8'b00000000; // d
		12'b01101111_1110: pixels <= 8'b00000000; // e
		12'b01101111_1111: pixels <= 8'b00000000; // f

		12'b01110000_0000: pixels <= 8'b00000000; // 0
		12'b01110000_0001: pixels <= 8'b00000000; // 1
		12'b01110000_0010: pixels <= 8'b00000000; // 2
		12'b01110000_0011: pixels <= 8'b00000000; // 3
		12'b01110000_0100: pixels <= 8'b00000000; // 4
		12'b01110000_0101: pixels <= 8'b11011100; // 5 ** ***
		12'b01110000_0110: pixels <= 8'b01100110; // 6  **  **
		12'b01110000_0111: pixels <= 8'b01100110; // 7  **  **
		12'b01110000_1000: pixels <= 8'b01100110; // 8  **  **
		12'b01110000_1001: pixels <= 8'b01100110; // 9  **  **
		12'b01110000_1010: pixels <= 8'b01100110; // a  **  **
		12'b01110000_1011: pixels <= 8'b01111100; // b  *****
		12'b01110000_1100: pixels <= 8'b01100000; // c  **
		12'b01110000_1101: pixels <= 8'b01100000; // d  **
		12'b01110000_1110: pixels <= 8'b11110000; // e ****
		12'b01110000_1111: pixels <= 8'b00000000; // f

		12'b01110001_0000: pixels <= 8'b00000000; // 0
		12'b01110001_0001: pixels <= 8'b00000000; // 1
		12'b01110001_0010: pixels <= 8'b00000000; // 2
		12'b01110001_0011: pixels <= 8'b00000000; // 3
		12'b01110001_0100: pixels <= 8'b00000000; // 4
		12'b01110001_0101: pixels <= 8'b01110110; // 5  *** **
		12'b01110001_0110: pixels <= 8'b11001100; // 6 **  **
		12'b01110001_0111: pixels <= 8'b11001100; // 7 **  **
		12'b01110001_1000: pixels <= 8'b11001100; // 8 **  **
		12'b01110001_1001: pixels <= 8'b11001100; // 9 **  **
		12'b01110001_1010: pixels <= 8'b11001100; // a **  **
		12'b01110001_1011: pixels <= 8'b01111100; // b  *****
		12'b01110001_1100: pixels <= 8'b00001100; // c     **
		12'b01110001_1101: pixels <= 8'b00001100; // d     **
		12'b01110001_1110: pixels <= 8'b00011110; // e    ****
		12'b01110001_1111: pixels <= 8'b00000000; // f

		12'b01110010_0000: pixels <= 8'b00000000; // 0
		12'b01110010_0001: pixels <= 8'b00000000; // 1
		12'b01110010_0010: pixels <= 8'b00000000; // 2
		12'b01110010_0011: pixels <= 8'b00000000; // 3
		12'b01110010_0100: pixels <= 8'b00000000; // 4
		12'b01110010_0101: pixels <= 8'b11011100; // 5 ** ***
		12'b01110010_0110: pixels <= 8'b01110110; // 6  *** **
		12'b01110010_0111: pixels <= 8'b01100110; // 7  **  **
		12'b01110010_1000: pixels <= 8'b01100000; // 8  **
		12'b01110010_1001: pixels <= 8'b01100000; // 9  **
		12'b01110010_1010: pixels <= 8'b01100000; // a  **
		12'b01110010_1011: pixels <= 8'b11110000; // b ****
		12'b01110010_1100: pixels <= 8'b00000000; // c
		12'b01110010_1101: pixels <= 8'b00000000; // d
		12'b01110010_1110: pixels <= 8'b00000000; // e
		12'b01110010_1111: pixels <= 8'b00000000; // f

		12'b01110011_0000: pixels <= 8'b00000000; // 0
		12'b01110011_0001: pixels <= 8'b00000000; // 1
		12'b01110011_0010: pixels <= 8'b00000000; // 2
		12'b01110011_0011: pixels <= 8'b00000000; // 3
		12'b01110011_0100: pixels <= 8'b00000000; // 4
		12'b01110011_0101: pixels <= 8'b01111100; // 5  *****
		12'b01110011_0110: pixels <= 8'b11000110; // 6 **   **
		12'b01110011_0111: pixels <= 8'b01100000; // 7  **
		12'b01110011_1000: pixels <= 8'b00111000; // 8   ***
		12'b01110011_1001: pixels <= 8'b00001100; // 9     **
		12'b01110011_1010: pixels <= 8'b11000110; // a **   **
		12'b01110011_1011: pixels <= 8'b01111100; // b  *****
		12'b01110011_1100: pixels <= 8'b00000000; // c
		12'b01110011_1101: pixels <= 8'b00000000; // d
		12'b01110011_1110: pixels <= 8'b00000000; // e
		12'b01110011_1111: pixels <= 8'b00000000; // f

		12'b01110100_0000: pixels <= 8'b00000000; // 0
		12'b01110100_0001: pixels <= 8'b00000000; // 1
		12'b01110100_0010: pixels <= 8'b00010000; // 2    *
		12'b01110100_0011: pixels <= 8'b00110000; // 3   **
		12'b01110100_0100: pixels <= 8'b00110000; // 4   **
		12'b01110100_0101: pixels <= 8'b11111100; // 5 ******
		12'b01110100_0110: pixels <= 8'b00110000; // 6   **
		12'b01110100_0111: pixels <= 8'b00110000; // 7   **
		12'b01110100_1000: pixels <= 8'b00110000; // 8   **
		12'b01110100_1001: pixels <= 8'b00110000; // 9   **
		12'b01110100_1010: pixels <= 8'b00110110; // a   ** **
		12'b01110100_1011: pixels <= 8'b00011100; // b    ***
		12'b01110100_1100: pixels <= 8'b00000000; // c
		12'b01110100_1101: pixels <= 8'b00000000; // d
		12'b01110100_1110: pixels <= 8'b00000000; // e
		12'b01110100_1111: pixels <= 8'b00000000; // f

		12'b01110101_0000: pixels <= 8'b00000000; // 0
		12'b01110101_0001: pixels <= 8'b00000000; // 1
		12'b01110101_0010: pixels <= 8'b00000000; // 2
		12'b01110101_0011: pixels <= 8'b00000000; // 3
		12'b01110101_0100: pixels <= 8'b00000000; // 4
		12'b01110101_0101: pixels <= 8'b11001100; // 5 **  **
		12'b01110101_0110: pixels <= 8'b11001100; // 6 **  **
		12'b01110101_0111: pixels <= 8'b11001100; // 7 **  **
		12'b01110101_1000: pixels <= 8'b11001100; // 8 **  **
		12'b01110101_1001: pixels <= 8'b11001100; // 9 **  **
		12'b01110101_1010: pixels <= 8'b11001100; // a **  **
		12'b01110101_1011: pixels <= 8'b01110110; // b  *** **
		12'b01110101_1100: pixels <= 8'b00000000; // c
		12'b01110101_1101: pixels <= 8'b00000000; // d
		12'b01110101_1110: pixels <= 8'b00000000; // e
		12'b01110101_1111: pixels <= 8'b00000000; // f

		12'b01110110_0000: pixels <= 8'b00000000; // 0
		12'b01110110_0001: pixels <= 8'b00000000; // 1
		12'b01110110_0010: pixels <= 8'b00000000; // 2
		12'b01110110_0011: pixels <= 8'b00000000; // 3
		12'b01110110_0100: pixels <= 8'b00000000; // 4
		12'b01110110_0101: pixels <= 8'b11000011; // 5 **    **
		12'b01110110_0110: pixels <= 8'b11000011; // 6 **    **
		12'b01110110_0111: pixels <= 8'b11000011; // 7 **    **
		12'b01110110_1000: pixels <= 8'b11000011; // 8 **    **
		12'b01110110_1001: pixels <= 8'b01100110; // 9  **  **
		12'b01110110_1010: pixels <= 8'b00111100; // a   ****
		12'b01110110_1011: pixels <= 8'b00011000; // b    **
		12'b01110110_1100: pixels <= 8'b00000000; // c
		12'b01110110_1101: pixels <= 8'b00000000; // d
		12'b01110110_1110: pixels <= 8'b00000000; // e
		12'b01110110_1111: pixels <= 8'b00000000; // f

		12'b01110111_0000: pixels <= 8'b00000000; // 0
		12'b01110111_0001: pixels <= 8'b00000000; // 1
		12'b01110111_0010: pixels <= 8'b00000000; // 2
		12'b01110111_0011: pixels <= 8'b00000000; // 3
		12'b01110111_0100: pixels <= 8'b00000000; // 4
		12'b01110111_0101: pixels <= 8'b11000011; // 5 **    **
		12'b01110111_0110: pixels <= 8'b11000011; // 6 **    **
		12'b01110111_0111: pixels <= 8'b11000011; // 7 **    **
		12'b01110111_1000: pixels <= 8'b11011011; // 8 ** ** **
		12'b01110111_1001: pixels <= 8'b11011011; // 9 ** ** **
		12'b01110111_1010: pixels <= 8'b11111111; // a ********
		12'b01110111_1011: pixels <= 8'b01100110; // b  **  **
		12'b01110111_1100: pixels <= 8'b00000000; // c
		12'b01110111_1101: pixels <= 8'b00000000; // d
		12'b01110111_1110: pixels <= 8'b00000000; // e
		12'b01110111_1111: pixels <= 8'b00000000; // f

		12'b01111000_0000: pixels <= 8'b00000000; // 0
		12'b01111000_0001: pixels <= 8'b00000000; // 1
		12'b01111000_0010: pixels <= 8'b00000000; // 2
		12'b01111000_0011: pixels <= 8'b00000000; // 3
		12'b01111000_0100: pixels <= 8'b00000000; // 4
		12'b01111000_0101: pixels <= 8'b11000011; // 5 **    **
		12'b01111000_0110: pixels <= 8'b01100110; // 6  **  **
		12'b01111000_0111: pixels <= 8'b00111100; // 7   ****
		12'b01111000_1000: pixels <= 8'b00011000; // 8    **
		12'b01111000_1001: pixels <= 8'b00111100; // 9   ****
		12'b01111000_1010: pixels <= 8'b01100110; // a  **  **
		12'b01111000_1011: pixels <= 8'b11000011; // b **    **
		12'b01111000_1100: pixels <= 8'b00000000; // c
		12'b01111000_1101: pixels <= 8'b00000000; // d
		12'b01111000_1110: pixels <= 8'b00000000; // e
		12'b01111000_1111: pixels <= 8'b00000000; // f

		12'b01111001_0000: pixels <= 8'b00000000; // 0
		12'b01111001_0001: pixels <= 8'b00000000; // 1
		12'b01111001_0010: pixels <= 8'b00000000; // 2
		12'b01111001_0011: pixels <= 8'b00000000; // 3
		12'b01111001_0100: pixels <= 8'b00000000; // 4
		12'b01111001_0101: pixels <= 8'b11000110; // 5 **   **
		12'b01111001_0110: pixels <= 8'b11000110; // 6 **   **
		12'b01111001_0111: pixels <= 8'b11000110; // 7 **   **
		12'b01111001_1000: pixels <= 8'b11000110; // 8 **   **
		12'b01111001_1001: pixels <= 8'b11000110; // 9 **   **
		12'b01111001_1010: pixels <= 8'b11000110; // a **   **
		12'b01111001_1011: pixels <= 8'b01111110; // b  ******
		12'b01111001_1100: pixels <= 8'b00000110; // c      **
		12'b01111001_1101: pixels <= 8'b00001100; // d     **
		12'b01111001_1110: pixels <= 8'b11111000; // e *****
		12'b01111001_1111: pixels <= 8'b00000000; // f

		12'b01111010_0000: pixels <= 8'b00000000; // 0
		12'b01111010_0001: pixels <= 8'b00000000; // 1
		12'b01111010_0010: pixels <= 8'b00000000; // 2
		12'b01111010_0011: pixels <= 8'b00000000; // 3
		12'b01111010_0100: pixels <= 8'b00000000; // 4
		12'b01111010_0101: pixels <= 8'b11111110; // 5 *******
		12'b01111010_0110: pixels <= 8'b11001100; // 6 **  **
		12'b01111010_0111: pixels <= 8'b00011000; // 7    **
		12'b01111010_1000: pixels <= 8'b00110000; // 8   **
		12'b01111010_1001: pixels <= 8'b01100000; // 9  **
		12'b01111010_1010: pixels <= 8'b11000110; // a **   **
		12'b01111010_1011: pixels <= 8'b11111110; // b *******
		12'b01111010_1100: pixels <= 8'b00000000; // c
		12'b01111010_1101: pixels <= 8'b00000000; // d
		12'b01111010_1110: pixels <= 8'b00000000; // e
		12'b01111010_1111: pixels <= 8'b00000000; // f

		default: pixels <= 8'b00000000;
    endcase
  end




endmodule
