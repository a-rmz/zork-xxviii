`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    23:57:42 05/10/2016
// Design Name:
// Module Name:    labyrynth_rom
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module labyrinth_rom(
    input [7:0] player_pos,
    input [7:0] screen_pos,
    output reg [7:0] char_ascii
    );

  always @ ( * ) begin
    case ( { player_pos, screen_pos } )


    // Position: (7, 7)
    16'b0111_0111_00000000: char_ascii = "A";
    16'b0111_0111_00000001: char_ascii = "l";
    16'b0111_0111_00000010: char_ascii = " ";
    16'b0111_0111_00000011: char_ascii = "o";
    16'b0111_0111_00000100: char_ascii = "e";
    16'b0111_0111_00000101: char_ascii = "s";
    16'b0111_0111_00000110: char_ascii = "t";
    16'b0111_0111_00000111: char_ascii = "e";
    16'b0111_0111_00001000: char_ascii = " ";
    16'b0111_0111_00001001: char_ascii = "s";
    16'b0111_0111_00001010: char_ascii = "e";
    16'b0111_0111_00001011: char_ascii = " ";
    16'b0111_0111_00001100: char_ascii = "i";
    16'b0111_0111_00001101: char_ascii = "m";
    16'b0111_0111_00001110: char_ascii = "p";
    16'b0111_0111_00001111: char_ascii = "o";
    16'b0111_0111_00010000: char_ascii = "n";
    16'b0111_0111_00010001: char_ascii = "e";
    16'b0111_0111_00010010: char_ascii = " ";
    16'b0111_0111_00010011: char_ascii = "u";
    16'b0111_0111_00010100: char_ascii = "n";
    16'b0111_0111_00010101: char_ascii = "a";
    16'b0111_0111_00010110: char_ascii = " ";
    16'b0111_0111_00010111: char_ascii = "g";
    16'b0111_0111_00011000: char_ascii = "r";
    16'b0111_0111_00011001: char_ascii = "a";
    16'b0111_0111_00011010: char_ascii = "n";
    16'b0111_0111_00011011: char_ascii = " ";
    16'b0111_0111_00011100: char_ascii = "m";
    16'b0111_0111_00011101: char_ascii = "o";
    16'b0111_0111_00011110: char_ascii = "n";
    16'b0111_0111_00011111: char_ascii = "t";
    16'b0111_0111_00100000: char_ascii = "a";
    16'b0111_0111_00100001: char_ascii = "n";
    16'b0111_0111_00100010: char_ascii = "a";
    16'b0111_0111_00100011: char_ascii = ".";
    16'b0111_0111_00100100: char_ascii = " ";
    16'b0111_0111_00100101: char_ascii = "N";
    16'b0111_0111_00100110: char_ascii = "o";
    16'b0111_0111_00100111: char_ascii = " ";
    16'b0111_0111_00101000: char_ascii = "e";
    16'b0111_0111_00101001: char_ascii = "r";
    16'b0111_0111_00101010: char_ascii = "e";
    16'b0111_0111_00101011: char_ascii = "s";
    16'b0111_0111_00101100: char_ascii = " ";
    16'b0111_0111_00101101: char_ascii = "c";
    16'b0111_0111_00101110: char_ascii = "a";
    16'b0111_0111_00101111: char_ascii = "p";
    16'b0111_0111_00110000: char_ascii = "a";
    16'b0111_0111_00110001: char_ascii = "z";
    16'b0111_0111_00110010: char_ascii = " ";
    16'b0111_0111_00110011: char_ascii = "d";
    16'b0111_0111_00110100: char_ascii = "e";
    16'b0111_0111_00110101: char_ascii = " ";
    16'b0111_0111_00110110: char_ascii = "d";
    16'b0111_0111_00110111: char_ascii = "i";
    16'b0111_0111_00111000: char_ascii = "s";
    16'b0111_0111_00111001: char_ascii = "t";
    16'b0111_0111_00111010: char_ascii = "i";
    16'b0111_0111_00111011: char_ascii = "n";
    16'b0111_0111_00111100: char_ascii = "g";
    16'b0111_0111_00111101: char_ascii = "u";
    16'b0111_0111_00111110: char_ascii = "i";
    16'b0111_0111_00111111: char_ascii = "r";
    16'b0111_0111_01000000: char_ascii = " ";
    16'b0111_0111_01000001: char_ascii = "n";
    16'b0111_0111_01000010: char_ascii = "a";
    16'b0111_0111_01000011: char_ascii = "d";
    16'b0111_0111_01000100: char_ascii = "a";
    16'b0111_0111_01000101: char_ascii = " ";
    16'b0111_0111_01000110: char_ascii = "s";
    16'b0111_0111_01000111: char_ascii = "a";
    16'b0111_0111_01001000: char_ascii = "l";
    16'b0111_0111_01001001: char_ascii = "v";
    16'b0111_0111_01001010: char_ascii = "o";
    16'b0111_0111_01001011: char_ascii = " ";
    16'b0111_0111_01001100: char_ascii = "p";
    16'b0111_0111_01001101: char_ascii = "r";
    16'b0111_0111_01001110: char_ascii = "o";
    16'b0111_0111_01001111: char_ascii = "f";
    16'b0111_0111_01010000: char_ascii = "u";
    16'b0111_0111_01010001: char_ascii = "n";
    16'b0111_0111_01010010: char_ascii = "d";
    16'b0111_0111_01010011: char_ascii = "a";
    16'b0111_0111_01010100: char_ascii = " ";
    16'b0111_0111_01010101: char_ascii = "o";
    16'b0111_0111_01010110: char_ascii = "s";
    16'b0111_0111_01010111: char_ascii = "c";
    16'b0111_0111_01011000: char_ascii = "u";
    16'b0111_0111_01011001: char_ascii = "r";
    16'b0111_0111_01011010: char_ascii = "i";
    16'b0111_0111_01011011: char_ascii = "d";
    16'b0111_0111_01011100: char_ascii = "a";
    16'b0111_0111_01011101: char_ascii = "d";
    16'b0111_0111_01011110: char_ascii = " ";
    16'b0111_0111_01011111: char_ascii = "e";
    16'b0111_0111_01100000: char_ascii = "n";
    16'b0111_0111_01100001: char_ascii = " ";
    16'b0111_0111_01100010: char_ascii = "l";
    16'b0111_0111_01100011: char_ascii = "a";
    16'b0111_0111_01100100: char_ascii = "s";
    16'b0111_0111_01100101: char_ascii = " ";
    16'b0111_0111_01100110: char_ascii = "d";
    16'b0111_0111_01100111: char_ascii = "e";
    16'b0111_0111_01101000: char_ascii = "m";
    16'b0111_0111_01101001: char_ascii = "a";
    16'b0111_0111_01101010: char_ascii = "s";
    16'b0111_0111_01101011: char_ascii = " ";
    16'b0111_0111_01101100: char_ascii = "d";
    16'b0111_0111_01101101: char_ascii = "i";
    16'b0111_0111_01101110: char_ascii = "r";
    16'b0111_0111_01101111: char_ascii = "e";
    16'b0111_0111_01110000: char_ascii = "c";
    16'b0111_0111_01110001: char_ascii = "c";
    16'b0111_0111_01110010: char_ascii = "i";
    16'b0111_0111_01110011: char_ascii = "o";
    16'b0111_0111_01110100: char_ascii = "n";
    16'b0111_0111_01110101: char_ascii = "e";
    16'b0111_0111_01110110: char_ascii = "s";
    16'b0111_0111_01110111: char_ascii = ".";
    16'b0111_0111_01111000: char_ascii = " ";
    16'b0111_0111_01111001: char_ascii = " ";
    16'b0111_0111_01111010: char_ascii = " ";
    16'b0111_0111_01111011: char_ascii = " ";
    16'b0111_0111_01111100: char_ascii = " ";
    16'b0111_0111_01111101: char_ascii = " ";
    16'b0111_0111_01111110: char_ascii = " ";
    16'b0111_0111_01111111: char_ascii = " ";
    16'b0111_0111_10000000: char_ascii = " ";
    16'b0111_0111_10000001: char_ascii = " ";
    16'b0111_0111_10000010: char_ascii = " ";
    16'b0111_0111_10000011: char_ascii = " ";
    16'b0111_0111_10000100: char_ascii = " ";
    16'b0111_0111_10000101: char_ascii = " ";
    16'b0111_0111_10000110: char_ascii = " ";
    16'b0111_0111_10000111: char_ascii = " ";
    16'b0111_0111_10001000: char_ascii = " ";
    16'b0111_0111_10001001: char_ascii = " ";
    16'b0111_0111_10001010: char_ascii = " ";
    16'b0111_0111_10001011: char_ascii = " ";
    16'b0111_0111_10001100: char_ascii = " ";
    16'b0111_0111_10001101: char_ascii = " ";
    16'b0111_0111_10001110: char_ascii = " ";
    16'b0111_0111_10001111: char_ascii = " ";
    16'b0111_0111_10010000: char_ascii = " ";
    16'b0111_0111_10010001: char_ascii = " ";
    16'b0111_0111_10010010: char_ascii = " ";
    16'b0111_0111_10010011: char_ascii = " ";
    16'b0111_0111_10010100: char_ascii = " ";
    16'b0111_0111_10010101: char_ascii = " ";
    16'b0111_0111_10010110: char_ascii = " ";
    16'b0111_0111_10010111: char_ascii = " ";
    16'b0111_0111_10011000: char_ascii = " ";
    16'b0111_0111_10011001: char_ascii = " ";
    16'b0111_0111_10011010: char_ascii = " ";
    16'b0111_0111_10011011: char_ascii = " ";
    16'b0111_0111_10011100: char_ascii = " ";
    16'b0111_0111_10011101: char_ascii = " ";
    16'b0111_0111_10011110: char_ascii = " ";
    16'b0111_0111_10011111: char_ascii = " ";
    16'b0111_0111_10100000: char_ascii = " ";
    16'b0111_0111_10100001: char_ascii = " ";
    16'b0111_0111_10100010: char_ascii = " ";
    16'b0111_0111_10100011: char_ascii = " ";
    16'b0111_0111_10100100: char_ascii = " ";
    16'b0111_0111_10100101: char_ascii = " ";
    16'b0111_0111_10100110: char_ascii = " ";
    16'b0111_0111_10100111: char_ascii = " ";
    16'b0111_0111_10101000: char_ascii = " ";
    16'b0111_0111_10101001: char_ascii = " ";
    16'b0111_0111_10101010: char_ascii = " ";
    16'b0111_0111_10101011: char_ascii = " ";
    16'b0111_0111_10101100: char_ascii = " ";
    16'b0111_0111_10101101: char_ascii = " ";
    16'b0111_0111_10101110: char_ascii = " ";
    16'b0111_0111_10101111: char_ascii = " ";
    16'b0111_0111_10110000: char_ascii = " ";
    16'b0111_0111_10110001: char_ascii = " ";
    16'b0111_0111_10110010: char_ascii = " ";
    16'b0111_0111_10110011: char_ascii = " ";
    16'b0111_0111_10110100: char_ascii = " ";
    16'b0111_0111_10110101: char_ascii = " ";
    16'b0111_0111_10110110: char_ascii = " ";
    16'b0111_0111_10110111: char_ascii = " ";
    16'b0111_0111_10111000: char_ascii = " ";
    16'b0111_0111_10111001: char_ascii = " ";
    16'b0111_0111_10111010: char_ascii = " ";
    16'b0111_0111_10111011: char_ascii = " ";
    16'b0111_0111_10111100: char_ascii = " ";
    16'b0111_0111_10111101: char_ascii = " ";
    16'b0111_0111_10111110: char_ascii = " ";
    16'b0111_0111_10111111: char_ascii = " ";
    16'b0111_0111_11000000: char_ascii = " ";
    16'b0111_0111_11000001: char_ascii = " ";
    16'b0111_0111_11000010: char_ascii = " ";
    16'b0111_0111_11000011: char_ascii = " ";
    16'b0111_0111_11000100: char_ascii = " ";
    16'b0111_0111_11000101: char_ascii = " ";
    16'b0111_0111_11000110: char_ascii = " ";
    16'b0111_0111_11000111: char_ascii = " ";
    16'b0111_0111_11001000: char_ascii = " ";
    16'b0111_0111_11001001: char_ascii = " ";
    16'b0111_0111_11001010: char_ascii = " ";
    16'b0111_0111_11001011: char_ascii = " ";
    16'b0111_0111_11001100: char_ascii = " ";
    16'b0111_0111_11001101: char_ascii = " ";
    16'b0111_0111_11001110: char_ascii = " ";
    16'b0111_0111_11001111: char_ascii = " ";
    16'b0111_0111_11010000: char_ascii = " ";
    16'b0111_0111_11010001: char_ascii = " ";
    16'b0111_0111_11010010: char_ascii = " ";
    16'b0111_0111_11010011: char_ascii = " ";
    16'b0111_0111_11010100: char_ascii = " ";
    16'b0111_0111_11010101: char_ascii = " ";
    16'b0111_0111_11010110: char_ascii = " ";
    16'b0111_0111_11010111: char_ascii = " ";
    16'b0111_0111_11011000: char_ascii = " ";
    16'b0111_0111_11011001: char_ascii = " ";
    16'b0111_0111_11011010: char_ascii = " ";
    16'b0111_0111_11011011: char_ascii = " ";
    16'b0111_0111_11011100: char_ascii = " ";
    16'b0111_0111_11011101: char_ascii = " ";
    16'b0111_0111_11011110: char_ascii = " ";
    16'b0111_0111_11011111: char_ascii = " ";
    16'b0111_0111_11100000: char_ascii = " ";
    16'b0111_0111_11100001: char_ascii = " ";
    16'b0111_0111_11100010: char_ascii = " ";
    16'b0111_0111_11100011: char_ascii = " ";
    16'b0111_0111_11100100: char_ascii = " ";
    16'b0111_0111_11100101: char_ascii = " ";
    16'b0111_0111_11100110: char_ascii = " ";
    16'b0111_0111_11100111: char_ascii = " ";
    16'b0111_0111_11101000: char_ascii = " ";
    16'b0111_0111_11101001: char_ascii = " ";
    16'b0111_0111_11101010: char_ascii = " ";
    16'b0111_0111_11101011: char_ascii = " ";
    16'b0111_0111_11101100: char_ascii = " ";
    16'b0111_0111_11101101: char_ascii = " ";
    16'b0111_0111_11101110: char_ascii = " ";
    16'b0111_0111_11101111: char_ascii = " ";
    16'b0111_0111_11110000: char_ascii = " ";
    16'b0111_0111_11110001: char_ascii = " ";
    16'b0111_0111_11110010: char_ascii = " ";
    16'b0111_0111_11110011: char_ascii = " ";
    16'b0111_0111_11110100: char_ascii = " ";
    16'b0111_0111_11110101: char_ascii = " ";
    16'b0111_0111_11110110: char_ascii = " ";
    16'b0111_0111_11110111: char_ascii = " ";
    16'b0111_0111_11111000: char_ascii = " ";
    16'b0111_0111_11111001: char_ascii = " ";
    16'b0111_0111_11111010: char_ascii = " ";
    16'b0111_0111_11111011: char_ascii = " ";
    16'b0111_0111_11111100: char_ascii = " ";
    16'b0111_0111_11111101: char_ascii = " ";
    16'b0111_0111_11111110: char_ascii = " ";
    16'b0111_0111_11111111: char_ascii = " ";

		default: char_ascii = " ";
    endcase
  end


endmodule
